`timescale 1ns/1ps

module inverter(input x, output y);
    assign y = ~x;
endmodule
