`timescale 1ns/1ps

module buf_gate(input x, output y);
    assign y = x;
endmodule
